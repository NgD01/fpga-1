//-----------------------------------------------------------------------------
//
// RAM image for input code file: hello.hex
//
//-----------------------------------------------------------------------------
module ram_image
(
	clk, addr, 
	we, din, dout
);
//-----------------------------------------------------------------------------
input           clk;
input   [11:0]  addr;
input           we;
input   [7:0]   din;
output  [7:0]   dout;
//-----------------------------------------------------------------------------
reg [7:0] dout;
reg [7:0] ram [4095:0];
//-----------------------------------------------------------------------------
initial 
begin
    ram[0] = 8'h21; ram[1] = 8'h00; ram[2] = 8'h0c; ram[3] = 8'hf9; 
    ram[4] = 8'hcd; ram[5] = 8'h30; ram[6] = 8'h03; ram[7] = 8'h00; 
    ram[8] = 8'hf5; ram[9] = 8'hc5; ram[10] = 8'hd5; ram[11] = 8'he5; 
    ram[12] = 8'hcd; ram[13] = 8'h24; ram[14] = 8'h03; ram[15] = 8'he1; 
    ram[16] = 8'hd1; ram[17] = 8'hc1; ram[18] = 8'hf1; ram[19] = 8'hfb; 
    ram[20] = 8'hc9; ram[21] = 8'h00; ram[22] = 8'h00; ram[23] = 8'h00; 
    ram[24] = 8'hf5; ram[25] = 8'hc5; ram[26] = 8'hd5; ram[27] = 8'he5; 
    ram[28] = 8'he1; ram[29] = 8'hd1; ram[30] = 8'hc1; ram[31] = 8'hf1; 
    ram[32] = 8'hfb; ram[33] = 8'hc9; ram[34] = 8'h00; ram[35] = 8'h00; 
    ram[36] = 8'h00; ram[37] = 8'h00; ram[38] = 8'h00; ram[39] = 8'h00; 
    ram[40] = 8'hf5; ram[41] = 8'hc5; ram[42] = 8'hd5; ram[43] = 8'he5; 
    ram[44] = 8'he1; ram[45] = 8'hd1; ram[46] = 8'hc1; ram[47] = 8'hf1; 
    ram[48] = 8'hfb; ram[49] = 8'hc9; ram[50] = 8'h00; ram[51] = 8'h00; 
    ram[52] = 8'h00; ram[53] = 8'h00; ram[54] = 8'h00; ram[55] = 8'h00; 
    ram[56] = 8'hf5; ram[57] = 8'hc5; ram[58] = 8'hd5; ram[59] = 8'he5; 
    ram[60] = 8'he1; ram[61] = 8'hd1; ram[62] = 8'hc1; ram[63] = 8'hf1; 
    ram[64] = 8'hfb; ram[65] = 8'hc9; ram[66] = 8'h7e; ram[67] = 8'h6f; 
    ram[68] = 8'h07; ram[69] = 8'h9f; ram[70] = 8'h67; ram[71] = 8'hc9; 
    ram[72] = 8'h7e; ram[73] = 8'h23; ram[74] = 8'h66; ram[75] = 8'h6f; 
    ram[76] = 8'hc9; ram[77] = 8'h7d; ram[78] = 8'h12; ram[79] = 8'hc9; 
    ram[80] = 8'h7d; ram[81] = 8'h12; ram[82] = 8'h13; ram[83] = 8'h7c; 
    ram[84] = 8'h12; ram[85] = 8'hc9; ram[86] = 8'h7d; ram[87] = 8'hb3; 
    ram[88] = 8'h6f; ram[89] = 8'h7c; ram[90] = 8'hb2; ram[91] = 8'h67; 
    ram[92] = 8'hc9; ram[93] = 8'h7d; ram[94] = 8'hab; ram[95] = 8'h6f; 
    ram[96] = 8'h7c; ram[97] = 8'haa; ram[98] = 8'h67; ram[99] = 8'hc9; 
    ram[100] = 8'h7d; ram[101] = 8'ha3; ram[102] = 8'h6f; ram[103] = 8'h7c; 
    ram[104] = 8'ha2; ram[105] = 8'h67; ram[106] = 8'hc9; ram[107] = 8'hcd; 
    ram[108] = 8'h91; ram[109] = 8'h00; ram[110] = 8'hc8; ram[111] = 8'h2b; 
    ram[112] = 8'hc9; ram[113] = 8'hcd; ram[114] = 8'h91; ram[115] = 8'h00; 
    ram[116] = 8'hc0; ram[117] = 8'h2b; ram[118] = 8'hc9; ram[119] = 8'heb; 
    ram[120] = 8'hcd; ram[121] = 8'h91; ram[122] = 8'h00; ram[123] = 8'hd8; 
    ram[124] = 8'h2b; ram[125] = 8'hc9; ram[126] = 8'hcd; ram[127] = 8'h91; 
    ram[128] = 8'h00; ram[129] = 8'hc8; ram[130] = 8'hd8; ram[131] = 8'h2b; 
    ram[132] = 8'hc9; ram[133] = 8'hcd; ram[134] = 8'h91; ram[135] = 8'h00; 
    ram[136] = 8'hd0; ram[137] = 8'h2b; ram[138] = 8'hc9; ram[139] = 8'hcd; 
    ram[140] = 8'h91; ram[141] = 8'h00; ram[142] = 8'hd8; ram[143] = 8'h2b; 
    ram[144] = 8'hc9; ram[145] = 8'h7b; ram[146] = 8'h95; ram[147] = 8'h5f; 
    ram[148] = 8'h7a; ram[149] = 8'h9c; ram[150] = 8'h21; ram[151] = 8'h01; 
    ram[152] = 8'h00; ram[153] = 8'hfa; ram[154] = 8'h9e; ram[155] = 8'h00; 
    ram[156] = 8'hb3; ram[157] = 8'hc9; ram[158] = 8'hb3; ram[159] = 8'h37; 
    ram[160] = 8'hc9; ram[161] = 8'hcd; ram[162] = 8'hbb; ram[163] = 8'h00; 
    ram[164] = 8'hd0; ram[165] = 8'h2b; ram[166] = 8'hc9; ram[167] = 8'hcd; 
    ram[168] = 8'hbb; ram[169] = 8'h00; ram[170] = 8'hd8; ram[171] = 8'h2b; 
    ram[172] = 8'hc9; ram[173] = 8'heb; ram[174] = 8'hcd; ram[175] = 8'hbb; 
    ram[176] = 8'h00; ram[177] = 8'hd8; ram[178] = 8'h2b; ram[179] = 8'hc9; 
    ram[180] = 8'hcd; ram[181] = 8'hbb; ram[182] = 8'h00; ram[183] = 8'hc8; 
    ram[184] = 8'hd8; ram[185] = 8'h2b; ram[186] = 8'hc9; ram[187] = 8'h7a; 
    ram[188] = 8'hbc; ram[189] = 8'hc2; ram[190] = 8'hc2; ram[191] = 8'h00; 
    ram[192] = 8'h7b; ram[193] = 8'hbd; ram[194] = 8'h21; ram[195] = 8'h01; 
    ram[196] = 8'h00; ram[197] = 8'hc9; ram[198] = 8'heb; ram[199] = 8'h7c; 
    ram[200] = 8'h17; ram[201] = 8'h7c; ram[202] = 8'h1f; ram[203] = 8'h67; 
    ram[204] = 8'h7d; ram[205] = 8'h1f; ram[206] = 8'h6f; ram[207] = 8'h1d; 
    ram[208] = 8'hc2; ram[209] = 8'hc7; ram[210] = 8'h00; ram[211] = 8'hc9; 
    ram[212] = 8'heb; ram[213] = 8'h29; ram[214] = 8'h1d; ram[215] = 8'hc2; 
    ram[216] = 8'hd5; ram[217] = 8'h00; ram[218] = 8'hc9; ram[219] = 8'h7b; 
    ram[220] = 8'h95; ram[221] = 8'h6f; ram[222] = 8'h7a; ram[223] = 8'h9c; 
    ram[224] = 8'h67; ram[225] = 8'hc9; ram[226] = 8'hcd; ram[227] = 8'he7; 
    ram[228] = 8'h00; ram[229] = 8'h23; ram[230] = 8'hc9; ram[231] = 8'h7c; 
    ram[232] = 8'h2f; ram[233] = 8'h67; ram[234] = 8'h7d; ram[235] = 8'h2f; 
    ram[236] = 8'h6f; ram[237] = 8'hc9; ram[238] = 8'h44; ram[239] = 8'h4d; 
    ram[240] = 8'h21; ram[241] = 8'h00; ram[242] = 8'h00; ram[243] = 8'h79; 
    ram[244] = 8'h0f; ram[245] = 8'hd2; ram[246] = 8'hf9; ram[247] = 8'h00; 
    ram[248] = 8'h19; ram[249] = 8'haf; ram[250] = 8'h78; ram[251] = 8'h1f; 
    ram[252] = 8'h47; ram[253] = 8'h79; ram[254] = 8'h1f; ram[255] = 8'h4f; 
    ram[256] = 8'hb0; ram[257] = 8'hc8; ram[258] = 8'haf; ram[259] = 8'h7b; 
    ram[260] = 8'h17; ram[261] = 8'h5f; ram[262] = 8'h7a; ram[263] = 8'h17; 
    ram[264] = 8'h57; ram[265] = 8'hb3; ram[266] = 8'hc8; ram[267] = 8'hc3; 
    ram[268] = 8'hf3; ram[269] = 8'h00; ram[270] = 8'h44; ram[271] = 8'h4d; 
    ram[272] = 8'h7a; ram[273] = 8'ha8; ram[274] = 8'hf5; ram[275] = 8'h7a; 
    ram[276] = 8'hb7; ram[277] = 8'hfc; ram[278] = 8'h4f; ram[279] = 8'h01; 
    ram[280] = 8'h78; ram[281] = 8'hb7; ram[282] = 8'hfc; ram[283] = 8'h57; 
    ram[284] = 8'h01; ram[285] = 8'h3e; ram[286] = 8'h10; ram[287] = 8'hf5; 
    ram[288] = 8'heb; ram[289] = 8'h11; ram[290] = 8'h00; ram[291] = 8'h00; 
    ram[292] = 8'h29; ram[293] = 8'hcd; ram[294] = 8'h5f; ram[295] = 8'h01; 
    ram[296] = 8'hca; ram[297] = 8'h3b; ram[298] = 8'h01; ram[299] = 8'hcd; 
    ram[300] = 8'h67; ram[301] = 8'h01; ram[302] = 8'hfa; ram[303] = 8'h3b; 
    ram[304] = 8'h01; ram[305] = 8'h7d; ram[306] = 8'hf6; ram[307] = 8'h01; 
    ram[308] = 8'h6f; ram[309] = 8'h7b; ram[310] = 8'h91; ram[311] = 8'h5f; 
    ram[312] = 8'h7a; ram[313] = 8'h98; ram[314] = 8'h57; ram[315] = 8'hf1; 
    ram[316] = 8'h3d; ram[317] = 8'hca; ram[318] = 8'h44; ram[319] = 8'h01; 
    ram[320] = 8'hf5; ram[321] = 8'hc3; ram[322] = 8'h24; ram[323] = 8'h01; 
    ram[324] = 8'hf1; ram[325] = 8'hf0; ram[326] = 8'hcd; ram[327] = 8'h4f; 
    ram[328] = 8'h01; ram[329] = 8'heb; ram[330] = 8'hcd; ram[331] = 8'h4f; 
    ram[332] = 8'h01; ram[333] = 8'heb; ram[334] = 8'hc9; ram[335] = 8'h7a; 
    ram[336] = 8'h2f; ram[337] = 8'h57; ram[338] = 8'h7b; ram[339] = 8'h2f; 
    ram[340] = 8'h5f; ram[341] = 8'h13; ram[342] = 8'hc9; ram[343] = 8'h78; 
    ram[344] = 8'h2f; ram[345] = 8'h47; ram[346] = 8'h79; ram[347] = 8'h2f; 
    ram[348] = 8'h4f; ram[349] = 8'h03; ram[350] = 8'hc9; ram[351] = 8'h7b; 
    ram[352] = 8'h17; ram[353] = 8'h5f; ram[354] = 8'h7a; ram[355] = 8'h17; 
    ram[356] = 8'h57; ram[357] = 8'hb3; ram[358] = 8'hc9; ram[359] = 8'h7b; 
    ram[360] = 8'h91; ram[361] = 8'h7a; ram[362] = 8'h98; ram[363] = 8'hc9; 
    ram[364] = 8'hdb; ram[365] = 8'h83; ram[366] = 8'hcd; ram[367] = 8'h43; 
    ram[368] = 8'h00; ram[369] = 8'he5; ram[370] = 8'h21; ram[371] = 8'h01; 
    ram[372] = 8'h00; ram[373] = 8'hd1; ram[374] = 8'hcd; ram[375] = 8'h64; 
    ram[376] = 8'h00; ram[377] = 8'h7c; ram[378] = 8'hb5; ram[379] = 8'hca; 
    ram[380] = 8'h81; ram[381] = 8'h01; ram[382] = 8'hc3; ram[383] = 8'h6c; 
    ram[384] = 8'h01; ram[385] = 8'h21; ram[386] = 8'h02; ram[387] = 8'h00; 
    ram[388] = 8'h39; ram[389] = 8'hcd; ram[390] = 8'h42; ram[391] = 8'h00; 
    ram[392] = 8'h7d; ram[393] = 8'hd3; ram[394] = 8'h80; ram[395] = 8'hc9; 
    ram[396] = 8'hdb; ram[397] = 8'h83; ram[398] = 8'hcd; ram[399] = 8'h43; 
    ram[400] = 8'h00; ram[401] = 8'he5; ram[402] = 8'h21; ram[403] = 8'h10; 
    ram[404] = 8'h00; ram[405] = 8'hd1; ram[406] = 8'hcd; ram[407] = 8'h64; 
    ram[408] = 8'h00; ram[409] = 8'h7c; ram[410] = 8'hb5; ram[411] = 8'hca; 
    ram[412] = 8'hae; ram[413] = 8'h01; ram[414] = 8'hdb; ram[415] = 8'h80; 
    ram[416] = 8'hcd; ram[417] = 8'h43; ram[418] = 8'h00; ram[419] = 8'h7d; 
    ram[420] = 8'h32; ram[421] = 8'h2c; ram[422] = 8'h04; ram[423] = 8'h21; 
    ram[424] = 8'h01; ram[425] = 8'h00; ram[426] = 8'hc9; ram[427] = 8'hc3; 
    ram[428] = 8'hb2; ram[429] = 8'h01; ram[430] = 8'h21; ram[431] = 8'h00; 
    ram[432] = 8'h00; ram[433] = 8'hc9; ram[434] = 8'hc9; ram[435] = 8'h21; 
    ram[436] = 8'h0d; ram[437] = 8'h00; ram[438] = 8'he5; ram[439] = 8'hcd; 
    ram[440] = 8'h6c; ram[441] = 8'h01; ram[442] = 8'hc1; ram[443] = 8'h21; 
    ram[444] = 8'h0a; ram[445] = 8'h00; ram[446] = 8'he5; ram[447] = 8'hcd; 
    ram[448] = 8'h6c; ram[449] = 8'h01; ram[450] = 8'hc1; ram[451] = 8'hc9; 
    ram[452] = 8'h21; ram[453] = 8'h02; ram[454] = 8'h00; ram[455] = 8'h39; 
    ram[456] = 8'hcd; ram[457] = 8'h48; ram[458] = 8'h00; ram[459] = 8'hcd; 
    ram[460] = 8'h42; ram[461] = 8'h00; ram[462] = 8'he5; ram[463] = 8'h21; 
    ram[464] = 8'h00; ram[465] = 8'h00; ram[466] = 8'hd1; ram[467] = 8'hcd; 
    ram[468] = 8'h71; ram[469] = 8'h00; ram[470] = 8'h7c; ram[471] = 8'hb5; 
    ram[472] = 8'hca; ram[473] = 8'hf4; ram[474] = 8'h01; ram[475] = 8'h21; 
    ram[476] = 8'h02; ram[477] = 8'h00; ram[478] = 8'h39; ram[479] = 8'he5; 
    ram[480] = 8'hcd; ram[481] = 8'h48; ram[482] = 8'h00; ram[483] = 8'h23; 
    ram[484] = 8'hd1; ram[485] = 8'hcd; ram[486] = 8'h50; ram[487] = 8'h00; 
    ram[488] = 8'h2b; ram[489] = 8'hcd; ram[490] = 8'h42; ram[491] = 8'h00; 
    ram[492] = 8'he5; ram[493] = 8'hcd; ram[494] = 8'h6c; ram[495] = 8'h01; 
    ram[496] = 8'hc1; ram[497] = 8'hc3; ram[498] = 8'hc4; ram[499] = 8'h01; 
    ram[500] = 8'hc9; ram[501] = 8'h21; ram[502] = 8'h02; ram[503] = 8'h00; 
    ram[504] = 8'h39; ram[505] = 8'hcd; ram[506] = 8'h48; ram[507] = 8'h00; 
    ram[508] = 8'he5; ram[509] = 8'h21; ram[510] = 8'h00; ram[511] = 8'h00; 
    ram[512] = 8'hd1; ram[513] = 8'hcd; ram[514] = 8'h8b; ram[515] = 8'h00; 
    ram[516] = 8'h7c; ram[517] = 8'hb5; ram[518] = 8'hca; ram[519] = 8'h24; 
    ram[520] = 8'h02; ram[521] = 8'h21; ram[522] = 8'h2d; ram[523] = 8'h00; 
    ram[524] = 8'he5; ram[525] = 8'hcd; ram[526] = 8'h6c; ram[527] = 8'h01; 
    ram[528] = 8'hc1; ram[529] = 8'h21; ram[530] = 8'h02; ram[531] = 8'h00; 
    ram[532] = 8'h39; ram[533] = 8'he5; ram[534] = 8'h21; ram[535] = 8'h04; 
    ram[536] = 8'h00; ram[537] = 8'h39; ram[538] = 8'hcd; ram[539] = 8'h48; 
    ram[540] = 8'h00; ram[541] = 8'hcd; ram[542] = 8'he2; ram[543] = 8'h00; 
    ram[544] = 8'hd1; ram[545] = 8'hcd; ram[546] = 8'h50; ram[547] = 8'h00; 
    ram[548] = 8'h21; ram[549] = 8'h02; ram[550] = 8'h00; ram[551] = 8'h39; 
    ram[552] = 8'hcd; ram[553] = 8'h48; ram[554] = 8'h00; ram[555] = 8'he5; 
    ram[556] = 8'hcd; ram[557] = 8'h31; ram[558] = 8'h02; ram[559] = 8'hc1; 
    ram[560] = 8'hc9; ram[561] = 8'hc5; ram[562] = 8'h21; ram[563] = 8'h00; 
    ram[564] = 8'h00; ram[565] = 8'h39; ram[566] = 8'he5; ram[567] = 8'h21; 
    ram[568] = 8'h06; ram[569] = 8'h00; ram[570] = 8'h39; ram[571] = 8'hcd; 
    ram[572] = 8'h48; ram[573] = 8'h00; ram[574] = 8'he5; ram[575] = 8'h21; 
    ram[576] = 8'h0a; ram[577] = 8'h00; ram[578] = 8'hd1; ram[579] = 8'hcd; 
    ram[580] = 8'h0e; ram[581] = 8'h01; ram[582] = 8'hd1; ram[583] = 8'hcd; 
    ram[584] = 8'h50; ram[585] = 8'h00; ram[586] = 8'h21; ram[587] = 8'h00; 
    ram[588] = 8'h00; ram[589] = 8'h39; ram[590] = 8'hcd; ram[591] = 8'h48; 
    ram[592] = 8'h00; ram[593] = 8'h7c; ram[594] = 8'hb5; ram[595] = 8'hca; 
    ram[596] = 8'h62; ram[597] = 8'h02; ram[598] = 8'h21; ram[599] = 8'h00; 
    ram[600] = 8'h00; ram[601] = 8'h39; ram[602] = 8'hcd; ram[603] = 8'h48; 
    ram[604] = 8'h00; ram[605] = 8'he5; ram[606] = 8'hcd; ram[607] = 8'h31; 
    ram[608] = 8'h02; ram[609] = 8'hc1; ram[610] = 8'h21; ram[611] = 8'h30; 
    ram[612] = 8'h00; ram[613] = 8'he5; ram[614] = 8'h21; ram[615] = 8'h06; 
    ram[616] = 8'h00; ram[617] = 8'h39; ram[618] = 8'hcd; ram[619] = 8'h48; 
    ram[620] = 8'h00; ram[621] = 8'he5; ram[622] = 8'h21; ram[623] = 8'h04; 
    ram[624] = 8'h00; ram[625] = 8'h39; ram[626] = 8'hcd; ram[627] = 8'h48; 
    ram[628] = 8'h00; ram[629] = 8'he5; ram[630] = 8'h21; ram[631] = 8'h0a; 
    ram[632] = 8'h00; ram[633] = 8'hd1; ram[634] = 8'hcd; ram[635] = 8'hee; 
    ram[636] = 8'h00; ram[637] = 8'hd1; ram[638] = 8'hcd; ram[639] = 8'hdb; 
    ram[640] = 8'h00; ram[641] = 8'hd1; ram[642] = 8'h19; ram[643] = 8'he5; 
    ram[644] = 8'hcd; ram[645] = 8'h6c; ram[646] = 8'h01; ram[647] = 8'hc1; 
    ram[648] = 8'hc1; ram[649] = 8'hc9; ram[650] = 8'hc5; ram[651] = 8'h21; 
    ram[652] = 8'h00; ram[653] = 8'h00; ram[654] = 8'h39; ram[655] = 8'he5; 
    ram[656] = 8'h21; ram[657] = 8'h06; ram[658] = 8'h00; ram[659] = 8'h39; 
    ram[660] = 8'hcd; ram[661] = 8'h48; ram[662] = 8'h00; ram[663] = 8'he5; 
    ram[664] = 8'h21; ram[665] = 8'h10; ram[666] = 8'h00; ram[667] = 8'hd1; 
    ram[668] = 8'hcd; ram[669] = 8'h0e; ram[670] = 8'h01; ram[671] = 8'hd1; 
    ram[672] = 8'hcd; ram[673] = 8'h50; ram[674] = 8'h00; ram[675] = 8'h21; 
    ram[676] = 8'h00; ram[677] = 8'h00; ram[678] = 8'h39; ram[679] = 8'hcd; 
    ram[680] = 8'h48; ram[681] = 8'h00; ram[682] = 8'h7c; ram[683] = 8'hb5; 
    ram[684] = 8'hca; ram[685] = 8'hbb; ram[686] = 8'h02; ram[687] = 8'h21; 
    ram[688] = 8'h00; ram[689] = 8'h00; ram[690] = 8'h39; ram[691] = 8'hcd; 
    ram[692] = 8'h48; ram[693] = 8'h00; ram[694] = 8'he5; ram[695] = 8'hcd; 
    ram[696] = 8'h8a; ram[697] = 8'h02; ram[698] = 8'hc1; ram[699] = 8'h21; 
    ram[700] = 8'h00; ram[701] = 8'h00; ram[702] = 8'h39; ram[703] = 8'he5; 
    ram[704] = 8'h21; ram[705] = 8'h06; ram[706] = 8'h00; ram[707] = 8'h39; 
    ram[708] = 8'hcd; ram[709] = 8'h48; ram[710] = 8'h00; ram[711] = 8'he5; 
    ram[712] = 8'h21; ram[713] = 8'h04; ram[714] = 8'h00; ram[715] = 8'h39; 
    ram[716] = 8'hcd; ram[717] = 8'h48; ram[718] = 8'h00; ram[719] = 8'he5; 
    ram[720] = 8'h21; ram[721] = 8'h10; ram[722] = 8'h00; ram[723] = 8'hd1; 
    ram[724] = 8'hcd; ram[725] = 8'hee; ram[726] = 8'h00; ram[727] = 8'hd1; 
    ram[728] = 8'hcd; ram[729] = 8'hdb; ram[730] = 8'h00; ram[731] = 8'hd1; 
    ram[732] = 8'hcd; ram[733] = 8'h50; ram[734] = 8'h00; ram[735] = 8'h21; 
    ram[736] = 8'h00; ram[737] = 8'h00; ram[738] = 8'h39; ram[739] = 8'hcd; 
    ram[740] = 8'h48; ram[741] = 8'h00; ram[742] = 8'he5; ram[743] = 8'h21; 
    ram[744] = 8'h09; ram[745] = 8'h00; ram[746] = 8'hd1; ram[747] = 8'hcd; 
    ram[748] = 8'h77; ram[749] = 8'h00; ram[750] = 8'h7c; ram[751] = 8'hb5; 
    ram[752] = 8'hca; ram[753] = 8'h10; ram[754] = 8'h03; ram[755] = 8'h21; 
    ram[756] = 8'h41; ram[757] = 8'h00; ram[758] = 8'he5; ram[759] = 8'h21; 
    ram[760] = 8'h02; ram[761] = 8'h00; ram[762] = 8'h39; ram[763] = 8'hcd; 
    ram[764] = 8'h48; ram[765] = 8'h00; ram[766] = 8'hd1; ram[767] = 8'h19; 
    ram[768] = 8'he5; ram[769] = 8'h21; ram[770] = 8'h0a; ram[771] = 8'h00; 
    ram[772] = 8'hd1; ram[773] = 8'hcd; ram[774] = 8'hdb; ram[775] = 8'h00; 
    ram[776] = 8'he5; ram[777] = 8'hcd; ram[778] = 8'h6c; ram[779] = 8'h01; 
    ram[780] = 8'hc1; ram[781] = 8'hc3; ram[782] = 8'h22; ram[783] = 8'h03; 
    ram[784] = 8'h21; ram[785] = 8'h30; ram[786] = 8'h00; ram[787] = 8'he5; 
    ram[788] = 8'h21; ram[789] = 8'h02; ram[790] = 8'h00; ram[791] = 8'h39; 
    ram[792] = 8'hcd; ram[793] = 8'h48; ram[794] = 8'h00; ram[795] = 8'hd1; 
    ram[796] = 8'h19; ram[797] = 8'he5; ram[798] = 8'hcd; ram[799] = 8'h6c; 
    ram[800] = 8'h01; ram[801] = 8'hc1; ram[802] = 8'hc1; ram[803] = 8'hc9; 
    ram[804] = 8'h21; ram[805] = 8'hd0; ram[806] = 8'h03; ram[807] = 8'he5; 
    ram[808] = 8'hcd; ram[809] = 8'hc4; ram[810] = 8'h01; ram[811] = 8'hc1; 
    ram[812] = 8'hcd; ram[813] = 8'hb3; ram[814] = 8'h01; ram[815] = 8'hc9; 
// jcw: change baud rate divisor from 195 to 163, for 19200 baud @ 50 MHz clock
//  ram[816] = 8'h21; ram[817] = 8'hc3; ram[818] = 8'h00; ram[819] = 8'h7d; 
    ram[816] = 8'h21; ram[817] = 8'ha3; ram[818] = 8'h00; ram[819] = 8'h7d; 
    ram[820] = 8'hd3; ram[821] = 8'h81; ram[822] = 8'h21; ram[823] = 8'h00; 
    ram[824] = 8'h00; ram[825] = 8'h7d; ram[826] = 8'hd3; ram[827] = 8'h82; 
    ram[828] = 8'h21; ram[829] = 8'h00; ram[830] = 8'h00; ram[831] = 8'h7d; 
    ram[832] = 8'hd3; ram[833] = 8'h84; ram[834] = 8'h21; ram[835] = 8'hff; 
    ram[836] = 8'h00; ram[837] = 8'h7d; ram[838] = 8'hd3; ram[839] = 8'h85; 
    ram[840] = 8'h21; ram[841] = 8'h00; ram[842] = 8'h00; ram[843] = 8'h7d; 
    ram[844] = 8'hd3; ram[845] = 8'h86; ram[846] = 8'h21; ram[847] = 8'hff; 
    ram[848] = 8'h00; ram[849] = 8'h7d; ram[850] = 8'hd3; ram[851] = 8'h87; 
    ram[852] = 8'h21; ram[853] = 8'h01; ram[854] = 8'h00; ram[855] = 8'h7d; 
    ram[856] = 8'hd3; ram[857] = 8'h88; ram[858] = 8'hfb; ram[859] = 8'h21; 
    ram[860] = 8'hea; ram[861] = 8'h03; ram[862] = 8'he5; ram[863] = 8'hcd; 
    ram[864] = 8'hc4; ram[865] = 8'h01; ram[866] = 8'hc1; ram[867] = 8'hcd; 
    ram[868] = 8'hb3; ram[869] = 8'h01; ram[870] = 8'h21; ram[871] = 8'hf9; 
    ram[872] = 8'h03; ram[873] = 8'he5; ram[874] = 8'hcd; ram[875] = 8'hc4; 
    ram[876] = 8'h01; ram[877] = 8'hc1; ram[878] = 8'h21; ram[879] = 8'h2d; 
    ram[880] = 8'h04; ram[881] = 8'he5; ram[882] = 8'h21; ram[883] = 8'h01; 
    ram[884] = 8'h00; ram[885] = 8'h29; ram[886] = 8'hd1; ram[887] = 8'h19; 
    ram[888] = 8'hcd; ram[889] = 8'h48; ram[890] = 8'h00; ram[891] = 8'he5; 
    ram[892] = 8'hcd; ram[893] = 8'hf5; ram[894] = 8'h01; ram[895] = 8'hc1; 
    ram[896] = 8'hcd; ram[897] = 8'hb3; ram[898] = 8'h01; ram[899] = 8'h21; 
    ram[900] = 8'h05; ram[901] = 8'h04; ram[902] = 8'he5; ram[903] = 8'hcd; 
    ram[904] = 8'hc4; ram[905] = 8'h01; ram[906] = 8'hc1; ram[907] = 8'h21; 
    ram[908] = 8'h2d; ram[909] = 8'h04; ram[910] = 8'he5; ram[911] = 8'h21; 
    ram[912] = 8'h00; ram[913] = 8'h00; ram[914] = 8'h29; ram[915] = 8'hd1; 
    ram[916] = 8'h19; ram[917] = 8'hcd; ram[918] = 8'h48; ram[919] = 8'h00; 
    ram[920] = 8'he5; ram[921] = 8'hcd; ram[922] = 8'h8a; ram[923] = 8'h02; 
    ram[924] = 8'hc1; ram[925] = 8'hcd; ram[926] = 8'hb3; ram[927] = 8'h01; 
    ram[928] = 8'h21; ram[929] = 8'h01; ram[930] = 8'h00; ram[931] = 8'h7d; 
    ram[932] = 8'hd3; ram[933] = 8'h84; ram[934] = 8'h21; ram[935] = 8'h13; 
    ram[936] = 8'h04; ram[937] = 8'he5; ram[938] = 8'hcd; ram[939] = 8'hc4; 
    ram[940] = 8'h01; ram[941] = 8'hc1; ram[942] = 8'hcd; ram[943] = 8'hb3; 
    ram[944] = 8'h01; ram[945] = 8'h21; ram[946] = 8'h01; ram[947] = 8'h00; 
    ram[948] = 8'h7c; ram[949] = 8'hb5; ram[950] = 8'hca; ram[951] = 8'hcf; 
    ram[952] = 8'h03; ram[953] = 8'hcd; ram[954] = 8'h8c; ram[955] = 8'h01; 
    ram[956] = 8'h7c; ram[957] = 8'hb5; ram[958] = 8'hca; ram[959] = 8'hcc; 
    ram[960] = 8'h03; ram[961] = 8'h3a; ram[962] = 8'h2c; ram[963] = 8'h04; 
    ram[964] = 8'hcd; ram[965] = 8'h43; ram[966] = 8'h00; ram[967] = 8'he5; 
    ram[968] = 8'hcd; ram[969] = 8'h6c; ram[970] = 8'h01; ram[971] = 8'hc1; 
    ram[972] = 8'hc3; ram[973] = 8'hb1; ram[974] = 8'h03; ram[975] = 8'hc9; 
    ram[976] = 8'h49; ram[977] = 8'h6e; ram[978] = 8'h74; ram[979] = 8'h65; 
    ram[980] = 8'h72; ram[981] = 8'h72; ram[982] = 8'h75; ram[983] = 8'h70; 
    ram[984] = 8'h74; ram[985] = 8'h20; ram[986] = 8'h30; ram[987] = 8'h20; 
    ram[988] = 8'h77; ram[989] = 8'h61; ram[990] = 8'h73; ram[991] = 8'h20; 
    ram[992] = 8'h61; ram[993] = 8'h73; ram[994] = 8'h73; ram[995] = 8'h65; 
    ram[996] = 8'h72; ram[997] = 8'h74; ram[998] = 8'h65; ram[999] = 8'h64; 
    ram[1000] = 8'h2e; ram[1001] = 8'h00; ram[1002] = 8'h48; ram[1003] = 8'h65; 
    ram[1004] = 8'h6c; ram[1005] = 8'h6c; ram[1006] = 8'h6f; ram[1007] = 8'h20; 
    ram[1008] = 8'h57; ram[1009] = 8'h6f; ram[1010] = 8'h72; ram[1011] = 8'h6c; 
    ram[1012] = 8'h64; ram[1013] = 8'h21; ram[1014] = 8'h21; ram[1015] = 8'h21; 
    ram[1016] = 8'h00; ram[1017] = 8'h44; ram[1018] = 8'h65; ram[1019] = 8'h63; 
    ram[1020] = 8'h20; ram[1021] = 8'h76; ram[1022] = 8'h61; ram[1023] = 8'h6c; 
    ram[1024] = 8'h75; ram[1025] = 8'h65; ram[1026] = 8'h3a; ram[1027] = 8'h20; 
    ram[1028] = 8'h00; ram[1029] = 8'h48; ram[1030] = 8'h65; ram[1031] = 8'h78; 
    ram[1032] = 8'h20; ram[1033] = 8'h76; ram[1034] = 8'h61; ram[1035] = 8'h6c; 
    ram[1036] = 8'h75; ram[1037] = 8'h65; ram[1038] = 8'h3a; ram[1039] = 8'h20; 
    ram[1040] = 8'h30; ram[1041] = 8'h78; ram[1042] = 8'h00; ram[1043] = 8'h45; 
    ram[1044] = 8'h63; ram[1045] = 8'h68; ram[1046] = 8'h6f; ram[1047] = 8'h69; 
    ram[1048] = 8'h6e; ram[1049] = 8'h67; ram[1050] = 8'h20; ram[1051] = 8'h72; 
    ram[1052] = 8'h65; ram[1053] = 8'h63; ram[1054] = 8'h65; ram[1055] = 8'h69; 
    ram[1056] = 8'h76; ram[1057] = 8'h65; ram[1058] = 8'h64; ram[1059] = 8'h20; 
    ram[1060] = 8'h62; ram[1061] = 8'h79; ram[1062] = 8'h74; ram[1063] = 8'h65; 
    ram[1064] = 8'h73; ram[1065] = 8'h3a; ram[1066] = 8'h20; ram[1067] = 8'h00; 
    ram[1068] = 8'h00; ram[1069] = 8'hd2; ram[1070] = 8'h04; ram[1071] = 8'h2e; 
    ram[1072] = 8'h16; ram[1073] = 8'h00; ram[1074] = 8'h00; ram[1075] = 8'h00; 
    ram[1076] = 8'h00; ram[1077] = 8'h00; ram[1078] = 8'h00; ram[1079] = 8'h00; 
    ram[1080] = 8'h00; ram[1081] = 8'h00; ram[1082] = 8'h00; ram[1083] = 8'h00; 
    ram[1084] = 8'h00; ram[1085] = 8'h00; ram[1086] = 8'h00; ram[1087] = 8'h00; 
    ram[1088] = 8'h00; ram[1089] = 8'h00; ram[1090] = 8'h00; ram[1091] = 8'h00; 
    ram[1092] = 8'h00; ram[1093] = 8'h00; ram[1094] = 8'h00; ram[1095] = 8'h00; 
    ram[1096] = 8'h00; ram[1097] = 8'h00; ram[1098] = 8'h00; ram[1099] = 8'h00; 
end

//-----------------------------------------------------------------------------
always @(posedge clk)
begin
    if (we)
    begin
        ram[addr] <= din;
        dout <= din;
    end
    else
        dout <= ram[addr];
end

endmodule
//-----------------------------------------------------------------------------
